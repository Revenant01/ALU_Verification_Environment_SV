package my_pkg;
  `include "Transaction.sv"
  `include "Generator.sv"
  `include "driver.sv"
  `include "Monitor.sv"
  `include "scoreboard.sv"
  `include "Environment.sv"
  `include "interface.sv"
  `include "test.sv"
  // `include "functional_Coverage.sv"
endpackage
